with address select
data <= 	x"00000021" when x"00000000",
	x"001b0006" when x"00000001",
	x"00020077" when x"00000002",
	x"fffd0037" when x"00000003",
	x"000006d0" when x"00000004",
	x"00000706" when x"00000005",
	x"0000e004" when x"00000006",
	x"00000036" when x"00000007",
	x"00040017" when x"00000008",
	x"00050077" when x"00000009",
	x"0001e706" when x"0000000a",
	x"fffb0037" when x"0000000b",
	x"000006d8" when x"0000000c",
	x"0000003b" when x"0000000d",
	x"000007d0" when x"0000000e",
	x"00050077" when x"0000000f",
	x"001a0784" when x"00000010",
	x"0000f00c" when x"00000011",
	x"000007d8" when x"00000012",
	x"0000003b" when x"00000013",
	x"00190784" when x"00000014",
	x"0000f744" when x"00000015",
	x"0001ef76" when x"00000016",
	x"fffe0017" when x"00000017",
	x"0000003b" when x"00000018",
	x"80000000" when x"00000019",
	x"80000001" when x"0000001a",
	x"00000048" when x"0000001b",
	x"00000065" when x"0000001c",
	x"0000006c" when x"0000001d",
	x"0000006c" when x"0000001e",
	x"0000006f" when x"0000001f",
	x"0000002c" when x"00000020",
	x"00000020" when x"00000021",
	x"00000057" when x"00000022",
	x"0000006f" when x"00000023",
	x"00000072" when x"00000024",
	x"0000006c" when x"00000025",
	x"00000064" when x"00000026",
	x"00000021" when x"00000027",
	x"00000000" when x"00000028",
	x"00000000" when others;
