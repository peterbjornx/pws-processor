clock_inst : clock PORT MAP (
		inclk	 => inclk_sig,
		outclk	 => outclk_sig
	);
